module test(
    input a, b,
    output out
);
    assign out = a & b; // Ví dụ đơn giản: AND hai tín hiệu
endmodule