`timescale 1ns/1ps
module fsqrt #(
    parameter WIDTH = 32
)(
    input   clk, rst_n, valid_input,
    input   [WIDTH-1:0] radicand,
    output  valid_output,
    output  [WIDTH-1:0] y
);
    reg [WIDTH-1:0] reg_a;
    wire [24:0]     f;
    wire [7:0]      res_e;
    wire [23:18]    Q23_18;
    wire [23:15]    Q23_15;
    wire [23:13]    Q23_13;
    wire [23:11]    Q23_11;
    wire [23:10]    Q23_10;
    wire [23:9]     Q23_9;
    wire [23:8]     Q23_8;
    wire [23:7]     Q23_7;
    wire [23:6]     Q23_6;
    wire [23:5]     Q23_5;
    wire [23:4]     Q23_4;
    wire [23:3]     Q23_3;
    wire [23:2]     Q23_2;
    wire [23:1]     Q23_1;
    wire [23:0]     Q23_0;

    wire [2:0]  A0, B0;
    wire [3:0]  X1, Y1, Z1, A1, B1;
    wire [4:0]  X2, Y2, Z2, A2, B2;
    wire [5:0]  X3, Y3, Z3, A3, B3;
    wire [6:0]  X4, Y4, Z4, A4, B4;
    wire [7:0]  X5, Y5, Z5, A5, B5;
    wire [8:0]  X6, Y6, Z6, A6, B6;
    wire [9:0]  X7, Y7, Z7, A7, B7;
    wire [10:0] X8, Y8, Z8, A8, B8;
    wire [11:0] X9, Y9, Z9, A9, B9;
    wire [12:0] X10, Y10, Z10, A10, B10;
    wire [13:0] X11, Y11, Z11, A11, B11;
    wire [14:0] X12, Y12, Z12, A12, B12;
    wire [15:0] X13, Y13, Z13, A13, B13;
    wire [16:0] X14, Y14, Z14, A14, B14;
    wire [17:0] X15, Y15, Z15, A15, B15;
    wire [18:0] X16, Y16, Z16, A16, B16;
    wire [19:0] X17, Y17, Z17, A17, B17;
    wire [20:0] X18, Y18, Z18, A18, B18;
    wire [21:0] X19, Y19, Z19, A19, B19;
    wire [22:0] X20, Y20, Z20, A20, B20;
    wire [23:0] X21, Y21, Z21, A21, B21;
    wire [24:0] X22, Y22, Z22, A22, B22;
    wire [25:0] X23, Y23, Z23, A23, B23;
    
    always @(posedge clk or negedge rst_n) begin
        if (~rst_n) begin
            reg_a <= 32'd0;
        end 
        else begin
            if(valid_input) begin
                reg_a <= radicand;
            end 
        end 
    end 

    reg         reg_s [0:13];
    reg [7:0]   reg_e [0:13];
    reg [12:0]  reg_f0;
    reg [6:0]   reg_f1;
    reg [2:0]   reg_f2;

    reg [7:0]   rsum0, rcar0;
    reg [10:0]  rsum1, rcar1;
    reg [12:0]  rsum2, rcar2;
    reg [14:0]  rsum3, rcar3;
    reg [15:0]  rsum4, rcar4;
    reg [16:0]  rsum5, rcar5;
    reg [17:0]  rsum6, rcar6;
    reg [18:0]  rsum7, rcar7;
    reg [19:0]  rsum8, rcar8;
    reg [20:0]  rsum9, rcar9;
    reg [21:0]  rsum10, rcar10;
    reg [22:0]  rsum11, rcar11;
    reg [23:0]  rsum12, rcar12;
    reg [24:0]  rsum13, rcar13;

    reg [5:0]   reg_Q23_18;
    reg [8:0]   reg_Q23_15;
    reg [10:0]  reg_Q23_13;
    reg [12:0]  reg_Q23_11;
    reg [13:0]  reg_Q23_10;
    reg [14:0]  reg_Q23_9;
    reg [15:0]  reg_Q23_8;
    reg [16:0]  reg_Q23_7;
    reg [17:0]  reg_Q23_6;
    reg [18:0]  reg_Q23_5;
    reg [19:0]  reg_Q23_4;
    reg [20:0]  reg_Q23_3;
    reg [21:0]  reg_Q23_2;
    reg [22:0]  reg_Q23_1;
    reg [23:0]  reg_Q23_0;
    reg [14:0]  reg_oValid;

    integer i;
    always @(posedge clk or negedge rst_n) begin
        if(~rst_n) begin
            for (i = 0; i < 14; i = i + 1'b1) begin
                reg_s[i] <= 1'b0;
                reg_e[i] <= 8'b0;
            end  
            reg_oValid  <= 15'd0;

            reg_f0  <= 13'd0;
            reg_f1  <= 7'd0;
            reg_f2  <= 3'd0;

            rsum0   <= 8'd0;
            rsum1   <= 11'd0;
            rsum2   <= 13'd0;
            rsum3   <= 15'd0;
            rsum4   <= 16'd0;
            rsum5   <= 17'd0;
            rsum6   <= 18'd0;
            rsum7   <= 19'd0;
            rsum8   <= 20'd0;
            rsum9   <= 21'd0;
            rsum10  <= 22'd0;
            rsum11  <= 23'd0;
            rsum12  <= 25'd0;
            rsum13  <= 25'd0;

            rcar0   <= 8'd0;
            rcar1   <= 11'd0;
            rcar2   <= 13'd0;
            rcar3   <= 15'd0;
            rcar4   <= 16'd0;
            rcar5   <= 17'd0;
            rcar6   <= 18'd0;
            rcar7   <= 19'd0;
            rcar8   <= 20'd0;
            rcar9   <= 21'd0;
            rcar10  <= 22'd0;
            rcar11  <= 23'd0;
            rcar12  <= 25'd0;
            rcar13  <= 25'd0;

            reg_Q23_18  <= 6'd0;
            reg_Q23_15  <= 9'd0; 
            reg_Q23_13  <= 11'd0;
            reg_Q23_11  <= 13'd0;
            reg_Q23_10  <= 14'd0;
            reg_Q23_9   <= 15'd0;
            reg_Q23_8   <= 16'd0;
            reg_Q23_7   <= 17'd0;
            reg_Q23_6   <= 18'd0;
            reg_Q23_5   <= 19'd0;
            reg_Q23_4   <= 20'd0;
            reg_Q23_3   <= 21'd0;
            reg_Q23_2   <= 22'd0;
            reg_Q23_1   <= 23'd0;
        end 
        else begin
            reg_oValid  <= {reg_oValid[13:0], valid_input};

            reg_s[0]    <= reg_a[31];
            reg_e[0]    <= res_e;
            reg_Q23_18  <= Q23_18;
            reg_f0      <= f[12:0];
            rsum0       <= A5;
            rcar0       <= B5;

            reg_s[1]    <= reg_s[0];
            reg_e[1]    <= reg_e[0];
            reg_Q23_15  <= Q23_15;
            reg_f1      <= reg_f0[6:0];
            rsum1       <= A8;
            rcar1       <= B8;

            reg_s[2]    <= reg_s[1];
            reg_e[2]    <= reg_e[1];
            reg_Q23_13  <= Q23_13;
            reg_f2      <= reg_f1[2:0];
            rsum2       <= A10;
            rcar2       <= B10;

            reg_s[3]    <= reg_s[2];
            reg_e[3]    <= reg_e[2];
            reg_Q23_11  <= Q23_11;
            rsum3       <= A12;
            rcar3       <= B12;

            reg_s[4]    <= reg_s[3];
            reg_e[4]    <= reg_e[3];
            reg_Q23_10  <= Q23_10;
            rsum4       <= A13;
            rcar4       <= B13;

            reg_s[5]    <= reg_s[4];
            reg_e[5]    <= reg_e[4];
            reg_Q23_9   <= Q23_9;
            rsum5       <= A14;
            rcar5       <= B14;

            reg_s[6]    <= reg_s[5];
            reg_e[6]    <= reg_e[5];
            reg_Q23_8   <= Q23_8;
            rsum6       <= A15;
            rcar6       <= B15;

            reg_s[7]    <= reg_s[6];
            reg_e[7]    <= reg_e[6];
            reg_Q23_7   <= Q23_7;
            rsum7       <= A16;
            rcar7       <= B16;

            reg_s[8]    <= reg_s[7];
            reg_e[8]    <= reg_e[7];
            reg_Q23_6   <= Q23_6;
            rsum8       <= A17;
            rcar8       <= B17;

            reg_s[9]    <= reg_s[8];
            reg_e[9]    <= reg_e[8];
            reg_Q23_5   <= Q23_5;
            rsum9       <= A18;
            rcar9       <= B18;

            reg_s[10]   <= reg_s[9];
            reg_e[10]   <= reg_e[9];
            reg_Q23_4   <= Q23_4;
            rsum10      <= A19;
            rcar10      <= B19;

            reg_s[11]   <= reg_s[10];
            reg_e[11]   <= reg_e[10];
            reg_Q23_3   <= Q23_3;
            rsum11      <= A20;
            rcar11      <= B20;

            reg_s[12]   <= reg_s[11];
            reg_e[12]   <= reg_e[11];
            reg_Q23_2   <= Q23_2;
            rsum12      <= A21;
            rcar12      <= B21;

            reg_s[13]   <= reg_s[12];
            reg_e[13]   <= reg_e[12];
            reg_Q23_1   <= Q23_1;
            rsum13      <= A22;
            rcar13      <= B22; 

            // reg_s[9]    <= reg_s[2];
            // reg_e[9]    <= reg_e[3];
            // reg_Q23_0  <= Q23_11;
        end 
    end 
    assign valid_output = reg_oValid[14];

    // ----------------------------------------- stage 1 -----------------------------------------
    assign res_e    = reg_a[30:24] + 8'd63 + reg_a[23];
    assign f        = (reg_a[23]) ? {2'b01, reg_a[22:0]} : {1'b1, reg_a[22:0], reg_a[0]};

    wire [3:0] T0       = {1'b0, A0} + {B0, 1'b0};
    assign Q23_18[23]   = ~T0[3];

    assign X1           = {A0[1:0], f[22:21]};
    assign Y1           = {Q23_18[23], 3'b011};
    assign Z1           = {B0[0], 3'b000};
    wire [4:0] T1       = {1'b0, A1} + {B1, 1'b0};
    assign Q23_18[22]   = ~T1[4];

    assign X2           = {A1[2:0], f[20:19]};
    assign Y2           = {Q23_18[22], Q23_18[22] ^ Q23_18[23], 3'b011};
    assign Z2           = {B1[1:0], 3'd0};
    wire [5:0] T2       = {1'b0, A2} + {B2, 1'b0};
    assign Q23_18[21]   = ~T2[5];

    assign X3           = {A2[3:0], f[18:17]};
    assign Y3           = {Q23_18[21], Q23_18[21] ^ Q23_18[22], Q23_18[21] ^ Q23_18[23], 3'b011};
    assign Z3           = {B2[2:0], 3'd0};
    wire [6:0] T3       = {1'b0, A3} + {B3, 1'b0};
    assign Q23_18[20]   = ~T3[6];

    assign X4           = {A3[4:0], f[16:15]};
    assign Y4           = {Q23_18[20], Q23_18[20] ^ Q23_18[23], Q23_18[20] ^ Q23_18[22], Q23_18[20] ^ Q23_18[21], 3'b011};
    assign Z4           = {B3[3:0], 3'd0};
    wire [7:0] T4       = {1'b0, A4} + {B4, 1'b0};
    assign Q23_18[19]   = ~T4[7];

    assign X5           = {A4[5:0], f[14:13]};
    assign Y5           = {Q23_18[19], Q23_18[19] ^ Q23_18[23], Q23_18[19] ^ Q23_18[22], Q23_18[19] ^ Q23_18[21],
                        Q23_18[19] ^ Q23_18[20], 3'b011};
    assign Z5           = {B4[4:0], 3'd0};
    wire [8:0] T5       = {1'b0, A5} + {B5, 1'b0};
    assign Q23_18[18]   = ~T5[8];


    // ----------------------------------------- stage 2 -----------------------------------------
    assign Q23_15[23:18]    = reg_Q23_18;
    assign X6               = {rsum0[6:0], reg_f0[12:11]};
    assign Y6               = {Q23_15[18],  Q23_15[18] ^ Q23_15[23], Q23_15[18] ^ Q23_15[22], Q23_15[18] ^ Q23_15[21], 
                                            Q23_15[18] ^ Q23_15[20], Q23_15[18] ^ Q23_15[19], 3'b011};
    assign Z6               = {rcar0[5:0], 3'd0};
    wire [9:0] T6           = {1'b0, A6} + {B6, 1'b0};
    assign Q23_15[17]       = ~T6[9];

    assign X7           = {A6[7:0], reg_f0[10:9]};
    assign Y7           = {Q23_15[17],  Q23_15[17] ^ Q23_15[23], Q23_15[17] ^ Q23_15[22], Q23_15[17] ^ Q23_15[21], Q23_15[17] ^ Q23_15[20], 
                                        Q23_15[17] ^ Q23_15[19], Q23_15[17] ^ Q23_15[18], 3'b011};
    assign Z7           = {B6[6:0], 3'd0};
    wire [10:0] T7      = {1'b0, A7} + {B7, 1'b0};
    assign Q23_15[16]   = ~T7[10];

    assign X8           = {A7[8:0], reg_f0[8:7]};
    assign Y8           = {Q23_15[16],  Q23_15[16] ^ Q23_15[23], Q23_15[16] ^ Q23_15[22], Q23_15[16] ^ Q23_15[21], Q23_15[16] ^ Q23_15[20], 
                                        Q23_15[16] ^ Q23_15[19], Q23_15[16] ^ Q23_15[18], Q23_15[16] ^ Q23_15[17], 3'b011};
    assign Z8           = {B7[7:0], 3'd0};
    wire [11:0] T8      = {1'b0, A8} + {B8, 1'b0};
    assign Q23_15[15]   = ~T8[11];

    // ----------------------------------------- stage 3 -----------------------------------------
    assign Q23_13[23:15] = reg_Q23_15;
    assign X9           = {rsum1[9:0], reg_f1[6:5]};
    assign Y9           = {Q23_13[15],  Q23_13[15] ^ Q23_13[23], Q23_13[15] ^ Q23_13[22], Q23_13[15] ^ Q23_13[21], 
                                        Q23_13[15] ^ Q23_13[20], Q23_13[15] ^ Q23_13[19], Q23_13[15] ^ Q23_13[18],
                                        Q23_13[15] ^ Q23_13[17], Q23_13[15] ^ Q23_13[16], 3'b011};
    assign Z9           = {rcar1[8:0], 3'd0};
    wire [12:0] T9      = {1'b0, A9} + {B9, 1'b0};
    assign Q23_13[14]   = ~T9[12];

    assign X10          = {A9[10:0], reg_f1[4:3]};
    assign Y10          = {Q23_13[14],  Q23_13[14] ^ Q23_13[23], Q23_13[14] ^ Q23_13[22], Q23_13[14] ^ Q23_13[21], 
                                        Q23_13[14] ^ Q23_13[20], Q23_13[14] ^ Q23_13[19], Q23_13[14] ^ Q23_13[18],
                                        Q23_13[14] ^ Q23_13[17], Q23_13[14] ^ Q23_13[16], Q23_13[14] ^ Q23_13[15], 3'b011};
    assign Z10          = {B9[9:0], 3'd0};
    wire [13:0] T10     = {1'b0, A10} + {B10, 1'b0};
    assign Q23_13[13]   = ~T10[13];

    // ----------------------------------------- stage 4 -----------------------------------------
    assign Q23_11[23:13] = reg_Q23_13;
    assign X11          = {rsum2[11:0], reg_f2[2:1]};
    assign Y11          = {Q23_11[13],  Q23_11[13] ^ Q23_11[23], Q23_11[13] ^ Q23_11[22], Q23_11[13] ^ Q23_11[21], 
                                        Q23_11[13] ^ Q23_11[20], Q23_11[13] ^ Q23_11[19], Q23_11[13] ^ Q23_11[18],
                                        Q23_11[13] ^ Q23_11[17], Q23_11[13] ^ Q23_11[16], Q23_11[13] ^ Q23_11[15], Q23_11[13] ^ Q23_11[14], 3'b011};
    assign Z11          = {rcar2[10:0], 3'd0};
    wire [14:0] T11     = {1'b0, A11} + {B11, 1'b0};
    assign Q23_11[12]   = ~T11[14];

    assign X12          = {A11[12:0], reg_f2[0], 1'b0};
    assign Y12          = {Q23_11[12],  Q23_11[12] ^ Q23_11[23], Q23_11[12] ^ Q23_11[22], Q23_11[12] ^ Q23_11[21], 
                                        Q23_11[12] ^ Q23_11[20], Q23_11[12] ^ Q23_11[19], Q23_11[12] ^ Q23_11[18],
                                        Q23_11[12] ^ Q23_11[17], Q23_11[12] ^ Q23_11[16], Q23_11[12] ^ Q23_11[15], 
                                        Q23_11[12] ^ Q23_11[14], Q23_11[12] ^ Q23_11[13], 3'b011};
    assign Z12          = {B11[11:0], 3'd0};
    wire [15:0] T12     = {1'b0, A12} + {B12, 1'b0};
    assign Q23_11[11]   = ~T12[15];

    // ----------------------------------------- stage 5 -----------------------------------------
    assign Q23_10[23:11] = reg_Q23_11;
    assign X13          = {rsum3[13:0], 2'b0};
    assign Y13          = {Q23_10[11],  Q23_10[11] ^ Q23_10[23], Q23_10[11] ^ Q23_10[22], Q23_10[11] ^ Q23_10[21], 
                                        Q23_10[11] ^ Q23_10[20], Q23_10[11] ^ Q23_10[19], Q23_10[11] ^ Q23_10[18],
                                        Q23_10[11] ^ Q23_10[17], Q23_10[11] ^ Q23_10[16], Q23_10[11] ^ Q23_10[15], 
                                        Q23_10[11] ^ Q23_10[14], Q23_10[11] ^ Q23_10[13], Q23_10[11] ^ Q23_10[12], 3'b011};
    assign Z13          = {rcar3[12:0], 3'd0};
    wire [16:0] T13     = {1'b0, A13} + {B13, 1'b0};
    assign Q23_10[10]   = ~T13[16];

    // ----------------------------------------- stage 6 -----------------------------------------
    assign Q23_9[23:10] = reg_Q23_10;
    assign X14          = {rsum4[14:0], 2'b0};
    assign Y14          = {Q23_9[10],   Q23_9[10] ^ Q23_9[23], Q23_9[10] ^ Q23_9[22], Q23_9[10] ^ Q23_9[21], 
                                        Q23_9[10] ^ Q23_9[20], Q23_9[10] ^ Q23_9[19], Q23_9[10] ^ Q23_9[18],
                                        Q23_9[10] ^ Q23_9[17], Q23_9[10] ^ Q23_9[16], Q23_9[10] ^ Q23_9[15], 
                                        Q23_9[10] ^ Q23_9[14], Q23_9[10] ^ Q23_9[13], Q23_9[10] ^ Q23_9[12],
                                        Q23_9[10] ^ Q23_9[11], 3'b011};
    assign Z14          = {rcar4[13:0], 3'd0};
    wire [17:0] T14     = {1'b0, A14} + {B14, 1'b0};
    assign Q23_9[9]     = ~T14[17];

    // ----------------------------------------- stage 7 -----------------------------------------
    assign Q23_8[23:9]  = reg_Q23_9;
    assign X15          = {rsum5[15:0], 2'b0};
    assign Y15          = {Q23_8[9],    Q23_8[9] ^ Q23_8[23], Q23_8[9] ^ Q23_8[22], Q23_8[9] ^ Q23_8[21], 
                                        Q23_8[9] ^ Q23_8[20], Q23_8[9] ^ Q23_8[19], Q23_8[9] ^ Q23_8[18],
                                        Q23_8[9] ^ Q23_8[17], Q23_8[9] ^ Q23_8[16], Q23_8[9] ^ Q23_8[15], 
                                        Q23_8[9] ^ Q23_8[14], Q23_8[9] ^ Q23_8[13], Q23_8[9] ^ Q23_8[12],
                                        Q23_8[9] ^ Q23_8[11], Q23_8[9] ^ Q23_8[10], 3'b011};
    assign Z15          = {rcar5[14:0], 3'd0};
    wire [18:0] T15     = {1'b0, A15} + {B15, 1'b0};
    assign Q23_8[8]     = ~T15[18];

    // ----------------------------------------- stage 8 -----------------------------------------
    assign Q23_7[23:8]  = reg_Q23_8;
    assign X16          = {rsum6[16:0], 2'b0};
    assign Y16          = {Q23_7[8],    Q23_7[8] ^ Q23_7[23], Q23_7[8] ^ Q23_7[22], Q23_7[8] ^ Q23_7[21], 
                                        Q23_7[8] ^ Q23_7[20], Q23_7[8] ^ Q23_7[19], Q23_7[8] ^ Q23_7[18],
                                        Q23_7[8] ^ Q23_7[17], Q23_7[8] ^ Q23_7[16], Q23_7[8] ^ Q23_7[15], 
                                        Q23_7[8] ^ Q23_7[14], Q23_7[8] ^ Q23_7[13], Q23_7[8] ^ Q23_7[12],
                                        Q23_7[8] ^ Q23_7[11], Q23_7[8] ^ Q23_7[10], Q23_7[8] ^ Q23_7[9], 3'b011};
    assign Z16          = {rcar6[15:0], 3'd0};
    wire [19:0] T16     = {1'b0, A16} + {B16, 1'b0};
    assign Q23_7[7]     = ~T16[19];

    // ----------------------------------------- stage 9 -----------------------------------------
    assign Q23_6[23:7]  = reg_Q23_7;
    assign X17          = {rsum7[17:0], 2'b0};
    assign Y17          = {Q23_6[7],    Q23_6[7] ^ Q23_6[23], Q23_6[7] ^ Q23_6[22], Q23_6[7] ^ Q23_6[21], 
                                        Q23_6[7] ^ Q23_6[20], Q23_6[7] ^ Q23_6[19], Q23_6[7] ^ Q23_6[18],
                                        Q23_6[7] ^ Q23_6[17], Q23_6[7] ^ Q23_6[16], Q23_6[7] ^ Q23_6[15], 
                                        Q23_6[7] ^ Q23_6[14], Q23_6[7] ^ Q23_6[13], Q23_6[7] ^ Q23_6[12],
                                        Q23_6[7] ^ Q23_6[11], Q23_6[7] ^ Q23_6[10], Q23_6[7] ^ Q23_6[9],
                                        Q23_6[7] ^ Q23_6[8] , 3'b011};
    assign Z17          = {rcar7[16:0], 3'd0};
    wire [20:0] T17     = {1'b0, A17} + {B17, 1'b0};
    assign Q23_6[6]     = ~T17[20];

    // ----------------------------------------- stage 10 -----------------------------------------
    assign Q23_5[23:6]  = reg_Q23_6;
    assign X18          = {rsum8[18:0], 2'b0};
    assign Y18          = {Q23_5[6],    Q23_5[6] ^ Q23_5[23], Q23_5[6] ^ Q23_5[22], Q23_5[6] ^ Q23_5[21], 
                                        Q23_5[6] ^ Q23_5[20], Q23_5[6] ^ Q23_5[19], Q23_5[6] ^ Q23_5[18],
                                        Q23_5[6] ^ Q23_5[17], Q23_5[6] ^ Q23_5[16], Q23_5[6] ^ Q23_5[15], 
                                        Q23_5[6] ^ Q23_5[14], Q23_5[6] ^ Q23_5[13], Q23_5[6] ^ Q23_5[12],
                                        Q23_5[6] ^ Q23_5[11], Q23_5[6] ^ Q23_5[10], Q23_5[6] ^ Q23_5[9],
                                        Q23_5[6] ^ Q23_5[8] , Q23_5[6] ^ Q23_5[7] , 3'b011};
    assign Z18          = {rcar8[17:0], 3'd0};
    wire [21:0] T18     = {1'b0, A18} + {B18, 1'b0};
    assign Q23_5[5]     = ~T18[21];

    // ----------------------------------------- stage 11 -----------------------------------------
    assign Q23_4[23:5]  = reg_Q23_5;
    assign X19          = {rsum9[19:0], 2'b0};
    assign Y19          = {Q23_4[5],    Q23_4[5] ^ Q23_4[23], Q23_4[5] ^ Q23_4[22], Q23_4[5] ^ Q23_4[21], 
                                        Q23_4[5] ^ Q23_4[20], Q23_4[5] ^ Q23_4[19], Q23_4[5] ^ Q23_4[18],
                                        Q23_4[5] ^ Q23_4[17], Q23_4[5] ^ Q23_4[16], Q23_4[5] ^ Q23_4[15], 
                                        Q23_4[5] ^ Q23_4[14], Q23_4[5] ^ Q23_4[13], Q23_4[5] ^ Q23_4[12],
                                        Q23_4[5] ^ Q23_4[11], Q23_4[5] ^ Q23_4[10], Q23_4[5] ^ Q23_4[9],
                                        Q23_4[5] ^ Q23_4[8] , Q23_4[5] ^ Q23_4[7] , Q23_4[5] ^ Q23_4[6], 3'b011};
    assign Z19          = {rcar9[18:0], 3'd0};
    wire [22:0] T19     = {1'b0, A19} + {B19, 1'b0};
    assign Q23_4[4]     = ~T19[22];

    // ----------------------------------------- stage 12 -----------------------------------------
    assign Q23_3[23:4]  = reg_Q23_4;
    assign X20          = {rsum10[20:0], 2'b0};
    assign Y20          = {Q23_3[4],    Q23_3[4] ^ Q23_3[23], Q23_3[4] ^ Q23_3[22], Q23_3[4] ^ Q23_3[21], 
                                        Q23_3[4] ^ Q23_3[20], Q23_3[4] ^ Q23_3[19], Q23_3[4] ^ Q23_3[18],
                                        Q23_3[4] ^ Q23_3[17], Q23_3[4] ^ Q23_3[16], Q23_3[4] ^ Q23_3[15], 
                                        Q23_3[4] ^ Q23_3[14], Q23_3[4] ^ Q23_3[13], Q23_3[4] ^ Q23_3[12],
                                        Q23_3[4] ^ Q23_3[11], Q23_3[4] ^ Q23_3[10], Q23_3[4] ^ Q23_3[9],
                                        Q23_3[4] ^ Q23_3[8] , Q23_3[4] ^ Q23_3[7] , Q23_3[4] ^ Q23_3[6],
                                        Q23_3[4] ^ Q23_3[5] , 3'b011};
    assign Z20          = {rcar10[19:0], 3'd0};
    wire [23:0] T20     = {1'b0, A20} + {B20, 1'b0};
    assign Q23_3[3]     = ~T20[23];

    // ----------------------------------------- stage 13 -----------------------------------------
    assign Q23_2[23:3]  = reg_Q23_3;
    assign X21          = {rsum11[21:0], 2'b0};
    assign Y21          = {Q23_2[3],    Q23_2[3] ^ Q23_2[23], Q23_2[3] ^ Q23_2[22], Q23_2[3] ^ Q23_2[21], 
                                        Q23_2[3] ^ Q23_2[20], Q23_2[3] ^ Q23_2[19], Q23_2[3] ^ Q23_2[18],
                                        Q23_2[3] ^ Q23_2[17], Q23_2[3] ^ Q23_2[16], Q23_2[3] ^ Q23_2[15], 
                                        Q23_2[3] ^ Q23_2[14], Q23_2[3] ^ Q23_2[13], Q23_2[3] ^ Q23_2[12],
                                        Q23_2[3] ^ Q23_2[11], Q23_2[3] ^ Q23_2[10], Q23_2[3] ^ Q23_2[9],
                                        Q23_2[3] ^ Q23_2[8] , Q23_2[3] ^ Q23_2[7] , Q23_2[3] ^ Q23_2[6],
                                        Q23_2[3] ^ Q23_2[5] , Q23_2[3] ^ Q23_2[4] , 3'b011};
    assign Z21          = {rcar11[20:0], 3'd0};
    wire [24:0] T21     = {1'b0, A21} + {B21, 1'b0};
    assign Q23_2[2]     = ~T21[24];

    // ----------------------------------------- stage 14 -----------------------------------------
    assign Q23_1[23:2]  = reg_Q23_2;
    assign X22          = {rsum12[22:0], 2'b0};
    assign Y22          = {Q23_2[2],    Q23_1[2] ^ Q23_1[23], Q23_1[2] ^ Q23_1[22], Q23_1[2] ^ Q23_1[21], 
                                        Q23_1[2] ^ Q23_1[20], Q23_1[2] ^ Q23_1[19], Q23_1[2] ^ Q23_1[18],
                                        Q23_1[2] ^ Q23_1[17], Q23_1[2] ^ Q23_1[16], Q23_1[2] ^ Q23_1[15], 
                                        Q23_1[2] ^ Q23_1[14], Q23_1[2] ^ Q23_1[13], Q23_1[2] ^ Q23_1[12],
                                        Q23_1[2] ^ Q23_1[11], Q23_1[2] ^ Q23_1[10], Q23_1[2] ^ Q23_1[9],
                                        Q23_1[2] ^ Q23_1[8] , Q23_1[2] ^ Q23_1[7] , Q23_1[2] ^ Q23_1[6],
                                        Q23_1[2] ^ Q23_1[5] , Q23_1[2] ^ Q23_1[4] , Q23_1[2] ^ Q23_1[3], 3'b011};
    assign Z22          = {rcar12[21:0], 3'd0};
    wire [25:0] T22     = {1'b0, A22} + {B22, 1'b0};
    assign Q23_1[1]     = ~T22[25];

    // ----------------------------------------- stage 15 -----------------------------------------
    assign Q23_0[23:1]  = reg_Q23_1;
    assign X23          = {rsum13[23:0], 2'b0};
    assign Y23          = {Q23_0[1],    Q23_0[1] ^ Q23_0[23], Q23_0[1] ^ Q23_0[22], Q23_0[1] ^ Q23_0[21], 
                                        Q23_0[1] ^ Q23_0[20], Q23_0[1] ^ Q23_0[19], Q23_0[1] ^ Q23_0[18],
                                        Q23_0[1] ^ Q23_0[17], Q23_0[1] ^ Q23_0[16], Q23_0[1] ^ Q23_0[15], 
                                        Q23_0[1] ^ Q23_0[14], Q23_0[1] ^ Q23_0[13], Q23_0[1] ^ Q23_0[12],
                                        Q23_0[1] ^ Q23_0[11], Q23_0[1] ^ Q23_0[10], Q23_0[1] ^ Q23_0[9],
                                        Q23_0[1] ^ Q23_0[8] , Q23_0[1] ^ Q23_0[7] , Q23_0[1] ^ Q23_0[6],
                                        Q23_0[1] ^ Q23_0[5] , Q23_0[1] ^ Q23_0[4] , Q23_0[1] ^ Q23_0[3],
                                        Q23_0[1] ^ Q23_0[2] , 3'b011};
    assign Z23          = {rcar13[22:0], 3'd0};
    wire [26:0] T23     = {1'b0, A23} + {B23, 1'b0};
    assign Q23_0[0]     = ~T23[26];

    assign y            = {reg_s[13], reg_e[13], Q23_0};

    csa #(.WIDTH(3))    csa0(.x({1'b0, f[24:23]}), .y(3'b111), .z(3'b000), .sum(A0), .carry(B0));
    csa #(.WIDTH(4))    csa1(.x(X1), .y(Y1), .z(Z1), .sum(A1), .carry(B1));
    csa #(.WIDTH(5))    csa2(.x(X2), .y(Y2), .z(Z2), .sum(A2), .carry(B2));
    csa #(.WIDTH(6))    csa3(.x(X3), .y(Y3), .z(Z3), .sum(A3), .carry(B3));
    csa #(.WIDTH(7))    csa4(.x(X4), .y(Y4), .z(Z4), .sum(A4), .carry(B4));
    csa #(.WIDTH(8))    csa5(.x(X5), .y(Y5), .z(Z5), .sum(A5), .carry(B5));

    csa #(.WIDTH(9))    csa6(.x(X6), .y(Y6), .z(Z6), .sum(A6), .carry(B6));
    csa #(.WIDTH(10))   csa7(.x(X7), .y(Y7), .z(Z7), .sum(A7), .carry(B7));
    csa #(.WIDTH(11))   csa8(.x(X8), .y(Y8), .z(Z8), .sum(A8), .carry(B8));

    csa #(.WIDTH(12))   csa9(.x(X9),   .y(Y9),  .z(Z9),  .sum(A9),  .carry(B9));
    csa #(.WIDTH(13))   csa10(.x(X10), .y(Y10), .z(Z10), .sum(A10), .carry(B10));

    csa #(.WIDTH(14))   csa11(.x(X11), .y(Y11), .z(Z11), .sum(A11), .carry(B11));
    csa #(.WIDTH(15))   csa12(.x(X12), .y(Y12), .z(Z12), .sum(A12), .carry(B12));

    csa #(.WIDTH(16))   csa13(.x(X13), .y(Y13), .z(Z13), .sum(A13), .carry(B13));
    csa #(.WIDTH(17))   csa14(.x(X14), .y(Y14), .z(Z14), .sum(A14), .carry(B14));
    csa #(.WIDTH(18))   csa15(.x(X15), .y(Y15), .z(Z15), .sum(A15), .carry(B15));
    csa #(.WIDTH(19))   csa16(.x(X16), .y(Y16), .z(Z16), .sum(A16), .carry(B16));
    csa #(.WIDTH(20))   csa17(.x(X17), .y(Y17), .z(Z17), .sum(A17), .carry(B17));
    csa #(.WIDTH(21))   csa18(.x(X18), .y(Y18), .z(Z18), .sum(A18), .carry(B18));
    csa #(.WIDTH(22))   csa19(.x(X19), .y(Y19), .z(Z19), .sum(A19), .carry(B19));
    csa #(.WIDTH(23))   csa20(.x(X20), .y(Y20), .z(Z20), .sum(A20), .carry(B20));
    csa #(.WIDTH(24))   csa21(.x(X21), .y(Y21), .z(Z21), .sum(A21), .carry(B21));
    csa #(.WIDTH(25))   csa22(.x(X22), .y(Y22), .z(Z22), .sum(A22), .carry(B22));
    csa #(.WIDTH(26))   csa23(.x(X23), .y(Y23), .z(Z23), .sum(A23), .carry(B23));
endmodule 