module RV32I();
endmodule