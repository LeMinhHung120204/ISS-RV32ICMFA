`timescale 1ns/1ps
module fsqrt2 #(
    parameter WIDTH = 32
)(
    input   clk, rst_n, valid_input,
    input   [WIDTH-1:0] radicand,
    output  valid_output,
    output  [WIDTH-1:0] y
);
    reg [WIDTH-1:0] reg_a;
    wire [24:0]     f;
    wire [7:0]      res_e;
    wire [23:18]    Q23_18;
    wire [23:15]    Q23_15;
    wire [23:13]    Q23_13;
    wire [23:11]    Q23_11;
    wire [23:10]    Q23_10;
    wire [23:9]     Q23_9;
    wire [23:8]     Q23_8;
    wire [23:7]     Q23_7;
    wire [23:6]     Q23_6;
    wire [23:5]     Q23_5;
    wire [23:4]     Q23_4;
    wire [23:3]     Q23_3;
    wire [23:2]     Q23_2;
    wire [23:1]     Q23_1;
    wire [23:0]     Q23_0;

    wire [2:0]  T0;
    wire [3:0]  T1;
    wire [4:0]  T2;
    wire [5:0]  T3; 
    wire [6:0]  T4;
    wire [7:0]  T5;
    wire [8:0]  A6, B6, C6, T6;
    wire [9:0]  A7, B7, C7, T7;
    wire [10:0] A8, B8, C8, T8;
    wire [11:0] A9, B9, C9, T9;
    wire [12:0] A10, B10, C10, T10;
    wire [13:0] A11, B11, C11, T11;
    wire [14:0] A12, B12, C12, T12;
    wire [15:0] A13, B13, C13, T13;
    wire [16:0] A14, B14, C14, T14;
    wire [17:0] A15, B15, C15, T15;
    wire [18:0] A16, B16, C16, T16;
    wire [19:0] A17, B17, C17, T17;
    wire [20:0] A18, B18, C18, T18;
    wire [21:0] A19, B19, C19, T19;
    wire [22:0] A20, B20, C20, T20;
    wire [23:0] A21, B21, C21, T21;
    wire [24:0] A22, B22, C22, T22;
    wire [25:0] A23, B23, C23, T23;
    
    always @(posedge clk or negedge rst_n) begin
        if (~rst_n) begin
            reg_a <= 32'd0;
        end 
        else begin
            if(valid_input) begin
                reg_a <= radicand;
            end 
        end 
    end 

    reg         reg_s [0:13];
    reg [7:0]   reg_e [0:13];
    reg [12:0]  reg_f0;
    reg [6:0]   reg_f1;
    reg [2:0]   reg_f2;

    reg [6:0]   rsum0;
    reg [9:0]   rsum1;
    reg [11:0]  rsum2;
    reg [13:0]  rsum3;
    reg [14:0]  rsum4;
    reg [15:0]  rsum5;
    reg [16:0]  rsum6;
    reg [17:0]  rsum7;
    reg [18:0]  rsum8;
    reg [19:0]  rsum9;
    reg [20:0]  rsum10;
    reg [21:0]  rsum11;
    reg [22:0]  rsum12;
    reg [23:0]  rsum13;

    reg [5:0]   reg_Q23_18;
    reg [8:0]   reg_Q23_15;
    reg [10:0]  reg_Q23_13;
    reg [12:0]  reg_Q23_11;
    reg [13:0]  reg_Q23_10;
    reg [14:0]  reg_Q23_9;
    reg [15:0]  reg_Q23_8;
    reg [16:0]  reg_Q23_7;
    reg [17:0]  reg_Q23_6;
    reg [18:0]  reg_Q23_5;
    reg [19:0]  reg_Q23_4;
    reg [20:0]  reg_Q23_3;
    reg [21:0]  reg_Q23_2;
    reg [22:0]  reg_Q23_1;
    reg [23:0]  reg_Q23_0;
    reg [14:0]  reg_oValid;

    integer i;
    always @(posedge clk or negedge rst_n) begin
        if(~rst_n) begin
            for (i = 0; i < 14; i = i + 1'b1) begin
                reg_s[i] <= 1'b0;
                reg_e[i] <= 8'b0;
            end  
            reg_oValid  <= 15'd0;

            reg_f0  <= 13'd0;
            reg_f1  <= 7'd0;
            reg_f2  <= 3'd0;

            rsum0   <= 7'd0;
            rsum1   <= 10'd0;
            rsum2   <= 12'd0;
            rsum3   <= 14'd0;
            rsum4   <= 15'd0;
            rsum5   <= 16'd0;
            rsum6   <= 17'd0;
            rsum7   <= 18'd0;
            rsum8   <= 19'd0;
            rsum9   <= 20'd0;
            rsum10  <= 21'd0;
            rsum11  <= 22'd0;
            rsum12  <= 23'd0;
            rsum13  <= 24'd0;

            reg_Q23_18  <= 6'd0;
            reg_Q23_15  <= 9'd0; 
            reg_Q23_13  <= 11'd0;
            reg_Q23_11  <= 13'd0;
            reg_Q23_10  <= 14'd0;
            reg_Q23_9   <= 15'd0;
            reg_Q23_8   <= 16'd0;
            reg_Q23_7   <= 17'd0;
            reg_Q23_6   <= 18'd0;
            reg_Q23_5   <= 19'd0;
            reg_Q23_4   <= 20'd0;
            reg_Q23_3   <= 21'd0;
            reg_Q23_2   <= 22'd0;
            reg_Q23_1   <= 23'd0;
        end 
        else begin
            reg_oValid  <= {reg_oValid[13:0], valid_input};
            rsum0       <= T5[6:0];
            reg_Q23_18  <= Q23_18;
            reg_e[0]    <= res_e;
            reg_f0      <= f[12:0];

            rsum1       <= T8[9:0];
            reg_Q23_15  <= Q23_15;
            reg_e[1]    <= reg_e[0];
            reg_f1      <= reg_f0[6:0];

            rsum2       <= T10[11:0];
            reg_Q23_13  <= Q23_13;
            reg_e[2]    <= reg_e[1];
            reg_f2      <= reg_f1[2:0];

            rsum3       <= T12[13:0];
            reg_Q23_11  <= Q23_11;
            reg_e[3]    <= reg_e[2];

            rsum4       <= T13[14:0];
            reg_Q23_10  <= Q23_10;
            reg_e[4]    <= reg_e[3];

            rsum5       <= T14[15:0];
            reg_Q23_9   <= Q23_9;
            reg_e[5]    <= reg_e[4];

            rsum6       <= T15[16:0];
            reg_Q23_8   <= Q23_8;
            reg_e[6]    <= reg_e[5];

            rsum7       <= T16[17:0];
            reg_Q23_7   <= Q23_7;
            reg_e[7]    <= reg_e[6];

            rsum8       <= T17[18:0];
            reg_Q23_6   <= Q23_6;
            reg_e[8]    <= reg_e[7];

            rsum9       <= T18[19:0];
            reg_Q23_5   <= Q23_5;
            reg_e[9]    <= reg_e[8];

            rsum10      <= T19[20:0];
            reg_Q23_4   <= Q23_4;
            reg_e[10]   <= reg_e[9];

            rsum11      <= T20[21:0];
            reg_Q23_3   <= Q23_3;
            reg_e[11]   <= reg_e[10];

            rsum12      <= T21[22:0];
            reg_Q23_2   <= Q23_2;
            reg_e[12]   <= reg_e[11];

            rsum13      <= T22[23:0];
            reg_Q23_1   <= Q23_1;
            reg_e[13]   <= reg_e[12];
        end 
    end 
    assign valid_output = reg_oValid[14];

    // ----------------------------------------- stage 1 -----------------------------------------
    assign res_e    = reg_a[30:24] + 8'd63 + reg_a[23];
    assign f        = (reg_a[23]) ? {2'b01, reg_a[22:0]} : {1'b1, reg_a[22:0], reg_a[0]};

    assign T0   = {1'b0, f[24:23]} - {3'b001};
    assign T1   = {T0[1:0], f[22:21]} + {~T0[2], 2'b01, T0[2]} + {3'b0, ~T0[2]};
    assign T2   = {T1[2:0], f[20:19]} + {~T1[3], T1[3] ^ T0[2], 2'b01, T1[3]} + {4'b0, ~T1[3]};
    assign T3   = {T2[3:0], f[18:17]} + {~T2[4], T2[4] ^ T0[2], T2[4] ^ T1[3], 2'b01, T2[4]} + {5'b0, ~T2[4]}; 
    assign T4   = {T3[4:0], f[16:15]} + {~T3[5], T3[5] ^ T0[2], T3[5] ^ T1[3], T3[5] ^ T2[4], 2'b01, T3[5]} + {6'b0, ~T3[5]};
    assign T5   = {T4[5:0], f[14:13]} + {~T4[6], T4[6] ^ T0[2], T4[6] ^ T1[3], T4[6] ^ T2[4], T4[6] ^ T3[5], 2'b01, T4[6]} + {7'b0, ~T4[6]};
    
    assign Q23_18[23] = ~T0[2];
    assign Q23_18[22] = ~T1[3];
    assign Q23_18[21] = ~T2[4];
    assign Q23_18[20] = ~T3[5];
    assign Q23_18[19] = ~T4[6];
    assign Q23_18[18] = ~T5[7];

    // ----------------------------------------- stage 1 -----------------------------------------
    assign Q23_15[23:18] = reg_Q23_18;
    assign A6 = {rsum0, reg_f0[12:11]};
    assign B6 = {Q23_15[18],    Q23_15[18] ^ Q23_15[23], Q23_15[18] ^ Q23_15[22], Q23_15[18] ^ Q23_15[21],
                                Q23_15[18] ^ Q23_15[20], Q23_15[18] ^ Q23_15[19], 2'b01, ~Q23_15[18]};
    assign C6 = {8'b0, Q23_15[18]};
    assign T6 = A6 + B6 + C6;
    assign Q23_15[17] = ~T6[8];

    assign A7 = {T6[7:0], reg_f0[10:9]};
    assign B7 = {Q23_15[17],    Q23_15[17] ^ Q23_15[23], Q23_15[17] ^ Q23_15[22], Q23_15[17] ^ Q23_15[21], 
                                Q23_15[17] ^ Q23_15[20], Q23_15[17] ^ Q23_15[19], Q23_15[17] ^ Q23_15[18], 2'b01, ~Q23_15[17]};
    assign C7 = {9'b0, Q23_15[17]};
    assign T7 = A7 + B7 + C7;
    assign Q23_15[16] = ~T7[9];

    assign A8 = {T7[8:0], reg_f0[8:7]};
    assign B8 = {Q23_15[16],    Q23_15[16] ^ Q23_15[23], Q23_15[16] ^ Q23_15[22], Q23_15[16] ^ Q23_15[21], Q23_15[16] ^ Q23_15[20], 
                                Q23_15[16] ^ Q23_15[19], Q23_15[16] ^ Q23_15[18], Q23_15[16] ^ Q23_15[17], 2'b01, ~Q23_15[16]};
    assign C8 = {10'b0, Q23_15[16]};
    assign T8 = A8 + B8 + C8;
    assign Q23_15[15] = ~T8[10];

    // ----------------------------------------- stage 2 -----------------------------------------
    wire [11:0] test = A9;

    assign Q23_13[23:15] = reg_Q23_15;
    assign A9 = {rsum1, reg_f1[6:5]};
    assign B9 = {Q23_13[15],    Q23_13[15] ^ Q23_13[23], Q23_13[15] ^ Q23_13[22], Q23_13[15] ^ Q23_13[21],
                                Q23_13[15] ^ Q23_13[20], Q23_13[15] ^ Q23_13[19], Q23_13[15] ^ Q23_13[18],
                                Q23_13[15] ^ Q23_13[17], Q23_13[15] ^ Q23_13[16], 2'b01, ~Q23_13[15]};
    assign C9 = Q23_13[15];
    assign T9 = A9 + B9 + C9;
    assign Q23_13[14] = ~T9[11];

    assign A10 = {T9[10:0], reg_f1[4:3]};
    assign B10 = {Q23_13[14],   Q23_13[14] ^ Q23_13[23], Q23_13[14] ^ Q23_13[22], Q23_13[14] ^ Q23_13[21], 
                                Q23_13[14] ^ Q23_13[20], Q23_13[14] ^ Q23_13[19], Q23_13[14] ^ Q23_13[18], 
                                Q23_13[14] ^ Q23_13[17], Q23_13[14] ^ Q23_13[16], Q23_13[14] ^ Q23_13[15], 2'b01, ~Q23_13[14]};
    assign C10 = Q23_13[14];
    assign T10 = A10 + B10 + C10;
    assign Q23_13[13] = ~T10[12];

    // ----------------------------------------- stage 3 -----------------------------------------
    assign Q23_11[23:13] = reg_Q23_13;
    assign A11 = {rsum2, reg_f2[2:1]};
    assign B11 = {Q23_11[13],   Q23_11[13] ^ Q23_11[23], Q23_11[13] ^ Q23_11[22], Q23_11[13] ^ Q23_11[21], 
                                Q23_11[13] ^ Q23_11[20], Q23_11[13] ^ Q23_11[19], Q23_11[13] ^ Q23_11[18], 
                                Q23_11[13] ^ Q23_11[17], Q23_11[13] ^ Q23_11[16], Q23_11[13] ^ Q23_11[15], 
                                Q23_11[13] ^ Q23_11[14], 2'b01, ~Q23_11[13]};
    assign C11 = Q23_11[13];
    assign T11 = A11 + B11 + C11;
    assign Q23_11[12] = ~T11[13];

    assign A12 = {T11[12:0], reg_f2[0], 1'b0};
    assign B12 = {Q23_11[12],   Q23_11[12] ^ Q23_11[23], Q23_11[12] ^ Q23_11[22], Q23_11[12] ^ Q23_11[21], 
                                Q23_11[12] ^ Q23_11[20], Q23_11[12] ^ Q23_11[19], Q23_11[12] ^ Q23_11[18], 
                                Q23_11[12] ^ Q23_11[17], Q23_11[12] ^ Q23_11[16], Q23_11[12] ^ Q23_11[15], 
                                Q23_11[12] ^ Q23_11[14], Q23_11[12] ^ Q23_11[13], 2'b01, ~Q23_11[12]};
    assign C12 = Q23_11[12];
    assign T12 = A12 + B12 + C12;
    assign Q23_11[11] = ~T12[14];

    // ----------------------------------------- stage 4 -----------------------------------------
    assign Q23_10[23:11] = reg_Q23_11;
    assign A13 = {rsum3, 2'b0};
    assign B13 = {Q23_10[11],   Q23_10[11] ^ Q23_10[23], Q23_10[11] ^ Q23_10[22], Q23_10[11] ^ Q23_10[21], 
                                Q23_10[11] ^ Q23_10[20], Q23_10[11] ^ Q23_10[19], Q23_10[11] ^ Q23_10[18], 
                                Q23_10[11] ^ Q23_10[17], Q23_10[11] ^ Q23_10[16], Q23_10[11] ^ Q23_10[15], 
                                Q23_10[11] ^ Q23_10[14], Q23_10[11] ^ Q23_10[13], Q23_10[11] ^ Q23_10[12], 2'b01,
                                ~Q23_10[11]};
    assign C13 = Q23_10[11];
    assign T13 = A13 + B13 + C13;
    assign Q23_10[10] = ~T13[15];

    // ----------------------------------------- stage 5 -----------------------------------------
    assign Q23_9[23:10] = reg_Q23_10;
    assign A14 = {rsum4, 2'b0};
    assign B14 = {Q23_9[10],    Q23_9[10] ^ Q23_9[23], Q23_9[10] ^ Q23_9[22], Q23_9[10] ^ Q23_9[21], 
                                Q23_9[10] ^ Q23_9[20], Q23_9[10] ^ Q23_9[19], Q23_9[10] ^ Q23_9[18], 
                                Q23_9[10] ^ Q23_9[17], Q23_9[10] ^ Q23_9[16], Q23_9[10] ^ Q23_9[15], 
                                Q23_9[10] ^ Q23_9[14], Q23_9[10] ^ Q23_9[13], Q23_9[10] ^ Q23_9[12], 
                                Q23_9[10] ^ Q23_9[11], 2'b01, ~Q23_9[10]};
    assign C14 = Q23_9[10];
    assign T14 = A14 + B14 + C14;
    assign Q23_9[9] = ~T14[16];

    // ----------------------------------------- stage 6 -----------------------------------------
    assign Q23_8[23:9] = reg_Q23_9;
    assign A15 = {rsum5, 2'b0};
    assign B15 = {Q23_8[9],     Q23_8[9] ^ Q23_8[23], Q23_8[9] ^ Q23_8[22], Q23_8[9] ^ Q23_8[21], 
                                Q23_8[9] ^ Q23_8[20], Q23_8[9] ^ Q23_8[19], Q23_8[9] ^ Q23_8[18], 
                                Q23_8[9] ^ Q23_8[17], Q23_8[9] ^ Q23_8[16], Q23_8[9] ^ Q23_8[15], 
                                Q23_8[9] ^ Q23_8[14], Q23_8[9] ^ Q23_8[13], Q23_8[9] ^ Q23_8[12], 
                                Q23_8[9] ^ Q23_8[11], Q23_8[9] ^ Q23_8[10], 2'b01, ~Q23_8[9]};
    assign C15 = Q23_8[9];
    assign T15 = A15 + B15 + C15;
    assign Q23_8[8] = ~T15[17];

    // ----------------------------------------- stage 7 -----------------------------------------
    assign Q23_7[23:8] = reg_Q23_8;
    assign A16 = {rsum6, 2'b0};
    assign B16 = {Q23_7[8], Q23_7[8] ^ Q23_7[23], Q23_7[8] ^ Q23_7[22], Q23_7[8] ^ Q23_7[21], 
                            Q23_7[8] ^ Q23_7[20], Q23_7[8] ^ Q23_7[19], Q23_7[8] ^ Q23_7[18], 
                            Q23_7[8] ^ Q23_7[17], Q23_7[8] ^ Q23_7[16], Q23_7[8] ^ Q23_7[15], 
                            Q23_7[8] ^ Q23_7[14], Q23_7[8] ^ Q23_7[13], Q23_7[8] ^ Q23_7[12], 
                            Q23_7[8] ^ Q23_7[11], Q23_7[8] ^ Q23_7[10], Q23_7[8] ^ Q23_7[9], 2'b01,
                            ~Q23_7[8]};
    assign C16 = Q23_7[8];
    assign T16 = A16 + B16 + C16;
    assign Q23_7[7] = ~T16[18];

    // ----------------------------------------- stage 8 -----------------------------------------
    assign Q23_6[23:7] = reg_Q23_7;
    assign A17 = {rsum7, 2'b0};
    assign B17 = {Q23_6[7], Q23_6[7] ^ Q23_6[23], Q23_6[7] ^ Q23_6[22], Q23_6[7] ^ Q23_6[21], 
                            Q23_6[7] ^ Q23_6[20], Q23_6[7] ^ Q23_6[19], Q23_6[7] ^ Q23_6[18], 
                            Q23_6[7] ^ Q23_6[17], Q23_6[7] ^ Q23_6[16], Q23_6[7] ^ Q23_6[15], 
                            Q23_6[7] ^ Q23_6[14], Q23_6[7] ^ Q23_6[13], Q23_6[7] ^ Q23_6[12], 
                            Q23_6[7] ^ Q23_6[11], Q23_6[7] ^ Q23_6[10], Q23_6[7] ^ Q23_6[9], 
                            Q23_6[7] ^ Q23_6[8] , 2'b01, ~Q23_6[7]};
    assign C17 = Q23_6[7];
    assign T17 = A17 + B17 + C17;
    assign Q23_6[6] = ~T17[19];
    
    // ----------------------------------------- stage 9 -----------------------------------------
    assign Q23_5[23:6] = reg_Q23_6;
    assign A18 = {rsum8, 2'b0};
    assign B18 = {Q23_5[6], Q23_5[6] ^ Q23_5[23], Q23_5[6] ^ Q23_5[22], Q23_5[6] ^ Q23_5[21], 
                            Q23_5[6] ^ Q23_5[20], Q23_5[6] ^ Q23_5[19], Q23_5[6] ^ Q23_5[18], 
                            Q23_5[6] ^ Q23_5[17], Q23_5[6] ^ Q23_5[16], Q23_5[6] ^ Q23_5[15], 
                            Q23_5[6] ^ Q23_5[14], Q23_5[6] ^ Q23_5[13], Q23_5[6] ^ Q23_5[12], 
                            Q23_5[6] ^ Q23_5[11], Q23_5[6] ^ Q23_5[10], Q23_5[6] ^ Q23_5[9], 
                            Q23_5[6] ^ Q23_5[8] , Q23_5[6] ^ Q23_5[7] , 2'b01, ~Q23_5[6]};
    assign C18 = Q23_5[6];
    assign T18 = A18 + B18 + C18;
    assign Q23_5[5] = ~T18[20];

    // ----------------------------------------- stage 10 -----------------------------------------
    assign Q23_4[23:5] = reg_Q23_5;
    assign A19 = {rsum9, 2'b0};
    assign B19 = {Q23_4[5], Q23_4[5] ^ Q23_4[23], Q23_4[5] ^ Q23_4[22], Q23_4[5] ^ Q23_4[21], 
                            Q23_4[5] ^ Q23_4[20], Q23_4[5] ^ Q23_4[19], Q23_4[5] ^ Q23_4[18], 
                            Q23_4[5] ^ Q23_4[17], Q23_4[5] ^ Q23_4[16], Q23_4[5] ^ Q23_4[15], 
                            Q23_4[5] ^ Q23_4[14], Q23_4[5] ^ Q23_4[13], Q23_4[5] ^ Q23_4[12], 
                            Q23_4[5] ^ Q23_4[11], Q23_4[5] ^ Q23_4[10], Q23_4[5] ^ Q23_4[9], 
                            Q23_4[5] ^ Q23_4[8] , Q23_4[5] ^ Q23_4[7] , Q23_4[5] ^ Q23_4[6], 
                            2'b01, ~Q23_4[5]};
    assign C19 = Q23_4[5];
    assign T19 = A19 + B19 + C19;
    assign Q23_4[4] = ~T19[21];

    // ----------------------------------------- stage 11 -----------------------------------------
    assign Q23_3[23:4] = reg_Q23_4;
    assign A20 = {rsum10, 2'b0};
    assign B20 = {Q23_3[4], Q23_3[4] ^ Q23_3[23], Q23_3[4] ^ Q23_3[22], Q23_3[4] ^ Q23_3[21], 
                            Q23_3[4] ^ Q23_3[20], Q23_3[4] ^ Q23_3[19], Q23_3[4] ^ Q23_3[18], 
                            Q23_3[4] ^ Q23_3[17], Q23_3[4] ^ Q23_3[16], Q23_3[4] ^ Q23_3[15], 
                            Q23_3[4] ^ Q23_3[14], Q23_3[4] ^ Q23_3[13], Q23_3[4] ^ Q23_3[12], 
                            Q23_3[4] ^ Q23_3[11], Q23_3[4] ^ Q23_3[10], Q23_3[4] ^ Q23_3[9], 
                            Q23_3[4] ^ Q23_3[8] , Q23_3[4] ^ Q23_3[7] , Q23_3[4] ^ Q23_3[6], 
                            Q23_3[4] ^ Q23_3[5] , 2'b01, ~Q23_3[4]};
    assign C20 = Q23_3[4];
    assign T20 = A20 + B20 + C20;
    assign Q23_3[3] = ~T20[22];

    // ----------------------------------------- stage 12 -----------------------------------------
    assign Q23_2[23:3] = reg_Q23_3;
    assign A21 = {rsum11, 2'b0};
    assign B21 = {Q23_2[3], Q23_2[3] ^ Q23_2[23], Q23_2[3] ^ Q23_2[22], Q23_2[3] ^ Q23_2[21], 
                            Q23_2[3] ^ Q23_2[20], Q23_2[3] ^ Q23_2[19], Q23_2[3] ^ Q23_2[18], 
                            Q23_2[3] ^ Q23_2[17], Q23_2[3] ^ Q23_2[15], Q23_2[3] ^ Q23_2[15], 
                            Q23_2[3] ^ Q23_2[14], Q23_2[3] ^ Q23_2[13], Q23_2[3] ^ Q23_2[12], 
                            Q23_2[3] ^ Q23_2[11], Q23_2[3] ^ Q23_2[10], Q23_2[3] ^ Q23_2[9], 
                            Q23_2[3] ^ Q23_2[8] , Q23_2[3] ^ Q23_2[7] , Q23_2[3] ^ Q23_2[6], 
                            Q23_2[3] ^ Q23_2[5] , Q23_2[3] ^ Q23_2[4] , 2'b01, ~Q23_2[3]};
    assign C21 = Q23_2[3];
    assign T21 = A21 + B21 + C21;
    assign Q23_2[2] = ~T21[23];

    // ----------------------------------------- stage 13 -----------------------------------------
    assign Q23_1[23:2] = reg_Q23_2;
    assign A22 = {rsum12, 2'b0};
    assign B22 = {Q23_1[2], Q23_1[2] ^ Q23_1[23], Q23_1[2] ^ Q23_1[22], Q23_1[2] ^ Q23_1[21], 
                            Q23_1[2] ^ Q23_1[20], Q23_1[2] ^ Q23_1[19], Q23_1[2] ^ Q23_1[18], 
                            Q23_1[2] ^ Q23_1[17], Q23_1[2] ^ Q23_1[16], Q23_1[2] ^ Q23_1[15], 
                            Q23_1[2] ^ Q23_1[14], Q23_1[2] ^ Q23_1[13], Q23_1[2] ^ Q23_1[12], 
                            Q23_1[2] ^ Q23_1[11], Q23_1[2] ^ Q23_1[10], Q23_1[2] ^ Q23_1[9], 
                            Q23_1[2] ^ Q23_1[8] , Q23_1[2] ^ Q23_1[7] , Q23_1[2] ^ Q23_1[6], 
                            Q23_1[2] ^ Q23_1[5] , Q23_1[2] ^ Q23_1[4] , Q23_1[2] ^ Q23_1[3], 
                            2'b01, ~Q23_1[2]};
    assign C22 = Q23_1[2];
    assign T22 = A22 + B22 + C22;
    assign Q23_1[1] = ~T22[24];

    // ----------------------------------------- stage 14 -----------------------------------------
    assign Q23_0[23:1] = reg_Q23_1;
    assign A23 = {rsum13, 2'b0};
    assign B23 = {Q23_0[1], Q23_0[1] ^ Q23_0[23], Q23_0[1] ^ Q23_0[22], Q23_0[1] ^ Q23_0[21], 
                            Q23_0[1] ^ Q23_0[20], Q23_0[1] ^ Q23_0[19], Q23_0[1] ^ Q23_0[18], 
                            Q23_0[1] ^ Q23_0[17], Q23_0[1] ^ Q23_0[16], Q23_0[1] ^ Q23_0[15], 
                            Q23_0[1] ^ Q23_0[14], Q23_0[1] ^ Q23_0[13], Q23_0[1] ^ Q23_0[12], 
                            Q23_0[1] ^ Q23_0[11], Q23_0[1] ^ Q23_0[10], Q23_0[1] ^ Q23_0[9], 
                            Q23_0[1] ^ Q23_0[8] , Q23_0[1] ^ Q23_0[7] , Q23_0[1] ^ Q23_0[6], 
                            Q23_0[1] ^ Q23_0[5] , Q23_0[1] ^ Q23_0[4] , Q23_0[1] ^ Q23_0[3], 
                            Q23_0[1] ^ Q23_0[2] , 2'b01, ~Q23_0[1]};
    assign C23 = Q23_0[1];
    assign T23 = A23 + B23 + C23;
    assign Q23_0[0] = ~T23[25];

    assign y = {1'b0, reg_e[13], Q23_0[22:0]};
    
endmodule 